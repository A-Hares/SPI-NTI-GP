`default_nettype none
`timescale 1ns/100ps

module SPI_TB;
    reg [7:0] SPCR_in

endmodule