`default_nettype none
module SCK_control(
    input wire M_BaudRate,
    input wire CPOL,
    input wire CPHA,
    output wire SCK_out,
    output wire Shift_clk,
    output wire Sample_clk
);


endmodule