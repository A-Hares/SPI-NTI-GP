//module top
